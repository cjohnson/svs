module tb;
  initial begin
    $display(0);
  end
endmodule
