module mux2to1(input logic test);
endmodule

