timeunit 100ps / 1fs;

module mux2to1(input logic test);
  timeunit 10ps; timeprecision 1fs;
endmodule

