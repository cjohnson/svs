module tb;
  initial begin
    $display("Hello world!");
    $display("This is a display statement!");
  end
endmodule
