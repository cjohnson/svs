module mux2to1(a[2:3] b[63:0]);
endmodule

module mux4to1();
endmodule
