module mux2to1;
endmodule

module mux4to1;
endmodule
