module tb;
  initial begin
    $display("");
  end
endmodule
