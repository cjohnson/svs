module tb;
  initial begin
    $display("Hello world!");
  end
endmodule
