module tb;
  initial begin
    $display("Hello world!\n");
  end
endmodule
