module mux2x1;
endmodule

