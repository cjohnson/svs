module m(output logic x);
  assign x = 2;
endmodule

module tb;
endmodule
