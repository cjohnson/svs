module tb;
  logic a;
  initial begin
    a = 1;
  end
endmodule
