module m(output logic x);
  assign x = 2;
endmodule

module tb;
  initial begin
    a = 2;
  end
endmodule
