module m(input logic x);
  assign x = 'h2;
endmodule
