timeunit 100ps / 1fs;

module mux2to1(input logic test);
endmodule

