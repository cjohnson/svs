module m(output logic x);
  assign x = 2;
endmodule

module tb;
  initial begin
    begin
    end
    begin end
  end
endmodule
